module CLA_4bit(a, b, cin, sum, cout);

endmodule


module CLA_4bit_P_G(a, b, cin, sum, P, G);

endmodule


module lookahead_carry_unit_16_bit(P0, G0, P1, G1, P2, G2, P3, G3, cin, C4, C8, C12, C16, GF, PF);

endmodule


module CLA_16bit(a, b, cin, sum, cout, Pout, Gout);

endmodule


module CLA_32bit(a, b, cin, sum, cout, Pout, Gout);

endmodule

module lookahead_carry_unit_32_bit (P0, G0, P1, G1, cin, C16, C32, GF, PF);

endmodule

