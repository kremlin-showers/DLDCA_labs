module half_adder(a, b, S, cout);

endmodule


module full_adder(a, b, cin, S, cout);

endmodule

module rca_Nbit #(parameter N = 32) (a, b, cin, S, cout);

endmodule


